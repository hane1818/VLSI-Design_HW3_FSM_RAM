entity My_ckt_3 is
port(
    clk, Read, Write: in bit;
    Data_Input: in bit_vector(7 downto 0);
    Data_Output: out bit_vector(7 downto 0));
end My_ckt_3;

architecture MODEL of My_ckt_3 is
begin

end MODEL;